library verilog;
use verilog.vl_types.all;
entity RAM_64bit_testbench is
end RAM_64bit_testbench;
