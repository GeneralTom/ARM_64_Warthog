module Program_Counter(out, in, PS, clock, reset);


	
	PC_DFF pc_dff ()
