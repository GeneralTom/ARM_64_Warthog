module GPIO_RM_testbench()
wire [63:0] data;
wire [15:0] IO;
wire [31:0] address;

reg [1:0] size;




endmodule
