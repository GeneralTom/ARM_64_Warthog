module PWM ();
    parameter base_address = 32'h80000000;

endmodule

module Timer_64 ();

endmodule

module Counter_64 (clock, reset, );
    input clock, reset
    
endmodule
