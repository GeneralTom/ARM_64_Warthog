// The branch logic goes in this file.
//
// You will need to look at both the ARM pdf, and
// The picture from the Discord.

module Branch_ControlUnit ();
	
endmodule
