module Datapath_With_Memory_testbench();
	
endmodule
