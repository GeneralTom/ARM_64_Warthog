// The data register logic goes in this file.
//
// You will need to look at both the ARM pdf, and
// The picture from the Discord.

module DataReg_ControlUnit ();

endmodule
