// The memory logic goes in this file.
//
// You will need to look at both the ARM pdf, and
// The picture from the Discord.

module Mem_ControlUnit ();

endmodule
